----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    17:09:00 04/10/2023 
-- Design Name: 
-- Module Name:    Decoder - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Decoder is
    Port ( Dec_IN : in  STD_LOGIC_VECTOR (4 downto 0);
           Dec_OUT : out  STD_LOGIC_VECTOR (31 downto 0));
end Decoder;

architecture Behavioral of Decoder is

begin

with Dec_IN select

	Dec_OUT <=  "0000_0000_0000_0000_0000_0000_0000_0001" when "00000",
					"0000_0000_0000_0000_0000_0000_0000_0010" when "00001",
					"0000_0000_0000_0000_0000_0000_0000_0100" when "00010",
					"0000_0000_0000_0000_0000_0000_0000_1000" when "00011",
					"0000_0000_0000_0000_0000_0000_0001_0000" when "00100",
					"0000_0000_0000_0000_0000_0000_0010_0000" when "00101",
					"0000_0000_0000_0000_0000_0000_0100_0000" when "00110",
					"0000_0000_0000_0000_0000_0000_1000_0000" when "00111",
					"0000_0000_0000_0000_0000_0001_0000_0000" when "01000",
					"0000_0000_0000_0000_0000_0010_0000_0000" when "01001",
					"0000_0000_0000_0000_0000_0100_0000_0000" when "01010",
					"0000_0000_0000_0000_0000_1000_0000_0000" when "01011",
					"0000_0000_0000_0000_0001_0000_0000_0000" when "01100",
					"0000_0000_0000_0000_0010_0000_0000_0000" when "01101",
					"0000_0000_0000_0000_0100_0000_0000_0000" when "01110",
					"0000_0000_0000_0000_1000_0000_0000_0000" when "01111",
					"0000_0000_0000_0001_0000_0000_0000_0000" when "10000",
					"0000_0000_0000_0010_0000_0000_0000_0000" when "10001",
					"0000_0000_0000_0100_0000_0000_0000_0000" when "10010",
					"0000_0000_0000_1000_0000_0000_0000_0000" when "10011",
					"0000_0000_0001_0000_0000_0000_0000_0000" when "10100",
					"0000_0000_0010_0000_0000_0000_0000_0000" when "10101",
					"0000_0000_0100_0000_0000_0000_0000_0000" when "10110",
					"0000_0000_1000_0000_0000_0000_0000_0000" when "10111",
					"0000_0001_0000_0000_0000_0000_0000_0000" when "11000",
					"0000_0010_0000_0000_0000_0000_0000_0000" when "11001",
					"0000_0100_0000_0000_0000_0000_0000_0000" when "11010",
					"0000_1000_0000_0000_0000_0000_0000_0000" when "11011",
					"0001_0000_0000_0000_0000_0000_0000_0000" when "11100",
					"0010_0000_0000_0000_0000_0000_0000_0000" when "11101",
					"0100_0000_0000_0000_0000_0000_0000_0000" when "11110",
					"1000_0000_0000_0000_0000_0000_0000_0000" when "11111",					

end Behavioral;

